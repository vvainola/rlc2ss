* Qucs 1.1.0 C:/Projects/rlc2ss/qucs/mutual_inductor.sch
.INCLUDE "C:/Programs/qucs_s_win64/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 1.1.0  C:/Projects/rlc2ss/qucs/mutual_inductor.sch
V1 _net0 0 DC 1
V2 _net1 0 DC 1
V3 _net2 0 DC 1
L1 _net3 _net6  1 
L2 _net4 _net6  1 
L3 _net5 _net6  1 
K12 L1 L2 0.9 
K21 L2 L3 0.9 
K31 L3 L1 0.9 
R1 _net0 _net3  10
R2 _net1 _net4  10
R3 _net2 _net5  10
VPr1 _net6 0 DC 0
.control
set filetype=ascii
op
print all > spice4qucs.cir.dc_op
destroy all
quit
.endc
.end
