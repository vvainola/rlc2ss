* Qucs 1.1.0 C:/Projects/rlc2ss/qucs/saturating_inductor.sch
.INCLUDE "C:/Programs/qucs_s_win64/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 1.1.0  C:/Projects/rlc2ss/qucs/saturating_inductor.sch
V _net0 0 DC 1
S1 _net0  _net2  _net3  _net4 
S2 _net2  _net5  _net6  _net7 
R 0 _net1  0.1
L0 _net1 _net0  0.01 
#DOUBLEL1=(0.015-0.01)/(2-1);
#DOUBLEL2=(0.0151-0.015)/(5-2);
#DOUBLEL1_ACT=(L1*L0)/(L0-L1);
#DOUBLEL2_ACT=(L2*L1_ACT)/(L1_ACT-L2);
L1 _net1 _net2  0.009999999999999997  IC=
L2 _net1 _net5  3.344481605351208E-5  IC=(0.0151-0.015)/(5-2)
.control
set filetype=ascii
op
print all > spice4qucs.cir.dc_op
destroy all
quit
.endc
.end
